

module rom_module (
    clk,
    address,
    q
    );
    
    input CLK;
    input [5:0]address;
    output [63:0]q;
    
    
    
endmodule

